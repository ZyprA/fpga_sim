module adder4(a,b,s);
    input [3:0] a, b;
    output [3:0] s;
    wire [2:0] c;

    assign s[0] = a[0] ^ b[0];
    assign c[0] = a[0] & b[0];
    assign s[1] = a[1] ^ b[1] ^ c[0];
    assign c[1] = (a[1] & b[1]) | (b[1] & c[0]) | (c[0] & a[1]);
    assign s[2] = a[2] ^ b[2] ^ c[1];
    assign c[2] = (a[2] & b[2]) | (b[2] & c[1]) | (c[1] & a[2]);
    assign s[3] = a[3] ^ b[3] ^ c[2];

endmodule

`timescale 1ns / 1ns

module adder4_sim;
    reg [3:0] a, b;
    wire [3:0] s;

    adder4 a4(a, b, s);

    initial begin
        $dumpfile("adder4.vcd");
        $dumpvars(0, adder4_sim);
    end

    initial begin
        a = 4'b0000; b = 4'b0000;
        #100 a = 4'b0001;
        #100 a = 4'b0010;
        #100 b = 4'b0111;
        #100 a = 4'b1101;
        #100 a = 4'b1011;
        #100 $finish;
    end

endmodule